module cpu(input wire clk, reset);
wire z,
     we3,
     wez,
     s_inc,
     selectorMuxSaltoR,
     selectorMuxRegistros,
     guardarMemoriaDatos,
     activarMemoriaDatos,
     selectorMuxDireccionesMemoriaDatos,
     activarPilaSubR,
     pushPilaSubR,
     selectorMuxPilaSubR,
     activarPilaDatos,
     pushPilaDatos,
     selectorMuxPilaDatos,
     selectorMuxAluMem_E_S;
wire [2:0] op_alu;
wire [5:0] opcode;

uc UnidadDeControl(opcode[5:0],
                   z,
                   clk,
                   we3,
                   wez,
                   s_inc,
                   selectorMuxSaltoR,
                   selectorMuxRegistros,
                   guardarMemoriaDatos,
                   activarMemoriaDatos,
                   selectorMuxDireccionesMemoriaDatos,
                   activarPilaSubR,
                   pushPilaSubR,
                   selectorMuxPilaSubR,
                   activarPilaDatos,
                   pushPilaDatos,
                   selectorMuxPilaDatos,
                   selectorMuxAluMem_E_S,
                   op_alu[2:0]);

cd CaminoDeDatos(clk,
                 reset,
                 we3,
                 wez,
                 s_inc,
                 selectorMuxSaltoR,
                 selectorMuxRegistros,
                 guardarMemoriaDatos,
                 activarMemoriaDatos,
                 selectorMuxDireccionesMemoriaDatos,
                 activarPilaSubR,
                 pushPilaSubR,
                 selectorMuxPilaSubR,
                 activarPilaDatos,
                 pushPilaDatos,
                 selectorMuxPilaDatos,
                 selectorMuxAluMem_E_S,
                 op_alu[2:0],
                 z,
                 opcode[5:0]);
endmodule
