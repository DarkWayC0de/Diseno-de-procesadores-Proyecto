module cpu(input wire clk, reset, 
   input wire [2:0] interrupciones,
           input wire [7:0] entradaDispositivo1,
           output wire [7:0] salidaDispositivo1,
           input wire [7:0] entradaDispositivo2,
           output wire [7:0] salidaDispositivo2,
           input wire [7:0] entradaDispositivo3,
           output wire [7:0] salidaDispositivo3,
           input wire [7:0] entradaDispositivo4,
           output wire [7:0] salidaDispositivo4,
           input wire [7:0] entradaDispositivo5,
           output wire [7:0] salidaDispositivo5);
wire z,
     we3,
     wez,
     s_inc,
     selectorMuxSaltoR,
     selectorMuxRegistros,
     guardarMemoriaDatos,
     activarMemoriaDatos,
     selectorMuxDireccionesMemoriaDatos,
     activarPilaSubR,
     pushPilaSubR,
     selectorMuxPilaSubR,
     activarPilaDatos,
     pushPilaDatos,
     selectorMuxPilaDatos,
     selectorMuxAluMem_E_S;
wire [2:0] op_alu;
wire [5:0] opcode;

uc UnidadDeControl(opcode[5:0],
                   z,
                   clk,
                   we3,
                   wez,
                   s_inc,
                   selectorMuxSaltoR,
                   selectorMuxRegistros,
                   guardarMemoriaDatos,
                   activarMemoriaDatos,
                   selectorMuxDireccionesMemoriaDatos,
                   activarPilaSubR,
                   pushPilaSubR,
                   selectorMuxPilaSubR,
                   activarPilaDatos,
                   pushPilaDatos,
                   selectorMuxPilaDatos,
                   selectorMuxAluMem_E_S,
                   op_alu[2:0]);

cd CaminoDeDatos(clk,
                 reset,
                 we3,
                 wez,
                 s_inc,
                 selectorMuxSaltoR,
                 selectorMuxRegistros,
                 guardarMemoriaDatos,
                 activarMemoriaDatos,
                 selectorMuxDireccionesMemoriaDatos,
                 activarPilaSubR,
                 pushPilaSubR,
                 selectorMuxPilaSubR,
                 activarPilaDatos,
                 pushPilaDatos,
                 selectorMuxPilaDatos,
                 selectorMuxAluMem_E_S,
                 op_alu[2:0],
                 interrupciones,
                 z,
                 opcode[5:0],
                 entradaDispositivo1 [7:0],
                 salidaDispositivo1 [7:0],
                 entradaDispositivo2 [7:0],
                 salidaDispositivo2 [7:0],
                 entradaDispositivo3 [7:0],
                 salidaDispositivo3 [7:0],
                 entradaDispositivo4 [7:0],
                 salidaDispositivo4 [7:0],
                 entradaDispositivo5 [7:0],
                 salidaDispositivo5 [7:0]);
endmodule
