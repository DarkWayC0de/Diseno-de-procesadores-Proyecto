module cpu(input wire clk, reset, 
           input wire [2:0] interrupciones,
	   output wire enable_whisbone,
           output wire rd, wr,
           output wire [15:0] dir,
           input wire [7:0] entradaDispositivo,
           output wire [7:0] salidaDispositivo);
wire z,
     we3,
     wez,
     s_inc,
     selectorMuxSaltoR,
     selectorMuxRegistros,
     guardarMemoriaDatos,
     activarMemoriaDatos,
     selectorMuxDireccionesMemoriaDatos,
     activarPilaSubR,
     pushPilaSubR,
     selectorMuxPilaSubR,
     activarPilaDatos,
     pushPilaDatos,
     selectorMuxPilaDatos,
     selectorMuxAluMem_E_S,
     editdirles,
     editdirhig;
wire [2:0] op_alu;
wire [5:0] opcode;

uc UnidadDeControl(opcode[5:0],
                   z,
                   clk,
                   we3,
                   wez,
                   s_inc,
                   selectorMuxSaltoR,
                   selectorMuxRegistros,
                   guardarMemoriaDatos,
                   activarMemoriaDatos,
                   selectorMuxDireccionesMemoriaDatos,
                   activarPilaSubR,
                   pushPilaSubR,
                   selectorMuxPilaSubR,
                   activarPilaDatos,
                   pushPilaDatos,
                   selectorMuxPilaDatos,
                   selectorMuxAluMem_E_S,
                   editdirles,
                   editdirhig,
                   op_alu[2:0]);

cd CaminoDeDatos(clk,
                 reset,
                 we3,
                 wez,
                 s_inc,
                 selectorMuxSaltoR,
                 selectorMuxRegistros,
                 guardarMemoriaDatos,
                 activarMemoriaDatos,
                 selectorMuxDireccionesMemoriaDatos,
                 activarPilaSubR,
                 pushPilaSubR,
                 selectorMuxPilaSubR,
                 activarPilaDatos,
                 pushPilaDatos,
                 selectorMuxPilaDatos,
                 selectorMuxAluMem_E_S,
                 editdirles,
                 editdirhig,
                 op_alu[2:0],
                 interrupciones,
                 z,
                 opcode[5:0],
                 rd, 
                 wr,
                 dir[15:0],
                 entradaDispositivo[7:0],
                 salidaDispositivo[7:0],
		 enable_wishbone
                 );
endmodule
