module cpu(input wire clk, reset);


endmodule
